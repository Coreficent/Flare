#version 400

in vec2 vertexPosition;
in vec4 vertexColor;
in vec2 vertexUV;

out vec2 fragmentPosition;
out vec4 fragmentColor;
out vec2 fragmentUV;

uniform mat4 cameraPosition;

void main() {
    gl_Position.xy = (cameraPosition * vec4(vertexPosition, 0.0, 1.0)).xy;
    gl_Position.z = 1.0;
    gl_Position.w = 1.0;
    
    fragmentPosition = vertexPosition;
    
    fragmentColor = vertexColor;
	
	fragmentUV = vec2(vertexUV.x, vertexUV.y);
}